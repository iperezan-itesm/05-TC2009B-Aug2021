/************************************************
  The Verilog HDL code example is from the book
  Computer Principles and Design in Verilog HDL
  by Yamin Li, published by A JOHN WILEY & SONS
************************************************/
module scinstmem_i2c_eeprom (a,inst); // instruction memory, rom
    input  [31:0] a;                  // address
    output [31:0] inst;               // instruction
    wire   [31:0] rom [0:127];        // rom cells: 128 words * 32 bits
    assign inst = rom[a[8:2]];        // use word address to read rom
    // rom[word_addr] = instruction
    assign rom[7'h00] = 32'b00110100000111010000000100000000;
    assign rom[7'h01] = 32'b00111100000010001100000000000000;
    assign rom[7'h02] = 32'b00111100000010011010000000000001;
    assign rom[7'h03] = 32'b00111100000000010000000000000000;
    assign rom[7'h04] = 32'b00110100001000010000000000000000;
    assign rom[7'h05] = 32'b00110100000001000000101001010101;
    assign rom[7'h06] = 32'b00110100000001110000000000000001;
    assign rom[7'h07] = 32'b10001100001001100000000000000000;
    assign rom[7'h08] = 32'b00000000000001100010111000000010;
    assign rom[7'h09] = 32'b00001100000000000000000000101011;
    assign rom[7'h0a] = 32'b00100000111001111111111111111111;
    assign rom[7'h0b] = 32'b00010000111000000000000000010101;
    assign rom[7'h0c] = 32'b00100000100001000000000000000001;
    assign rom[7'h0d] = 32'b00000000000001100010101000000000;
    assign rom[7'h0e] = 32'b00000000000001010010111000000010;
    assign rom[7'h0f] = 32'b00001100000000000000000000101011;
    assign rom[7'h10] = 32'b00100000111001111111111111111111;
    assign rom[7'h11] = 32'b00010000111000000000000000001111;
    assign rom[7'h12] = 32'b00100000100001000000000000000001;
    assign rom[7'h13] = 32'b00000000000001100010110000000000;
    assign rom[7'h14] = 32'b00000000000001010010111000000010;
    assign rom[7'h15] = 32'b00001100000000000000000000101011;
    assign rom[7'h16] = 32'b00100000111001111111111111111111;
    assign rom[7'h17] = 32'b00010000111000000000000000001001;
    assign rom[7'h18] = 32'b00100000100001000000000000000001;
    assign rom[7'h19] = 32'b00000000000001100010111000000000;
    assign rom[7'h1a] = 32'b00000000000001010010111000000010;
    assign rom[7'h1b] = 32'b00001100000000000000000000101011;
    assign rom[7'h1c] = 32'b00100000111001111111111111111111;
    assign rom[7'h1d] = 32'b00010000111000000000000000000011;
    assign rom[7'h1e] = 32'b00100000100001000000000000000001;
    assign rom[7'h1f] = 32'b00100000001000010000000000000100;
    assign rom[7'h20] = 32'b00001000000000000000000000000111;
    assign rom[7'h21] = 32'b00110100000001000000101001010101;
    assign rom[7'h22] = 32'b00110100000001110000000000000001;
    assign rom[7'h23] = 32'b00001100000000000000000000111001;
    assign rom[7'h24] = 32'b10101101000000100000000000000000;
    assign rom[7'h25] = 32'b00100001000010000000000000000100;
    assign rom[7'h26] = 32'b00100000100001000000000000000001;
    assign rom[7'h27] = 32'b00100000111001111111111111111111;
    assign rom[7'h28] = 32'b00010000111000000000000000000001;
    assign rom[7'h29] = 32'b00001000000000000000000000100011;
    assign rom[7'h2a] = 32'b00001000000000000000000000101010;
    assign rom[7'h2b] = 32'b00100011101111011111111111110000;
    assign rom[7'h2c] = 32'b10101111101111110000000000001100;
    assign rom[7'h2d] = 32'b10101111101111100000000000001000;
    assign rom[7'h2e] = 32'b00000000000111011111000000000000;
    assign rom[7'h2f] = 32'b00001100000000000000000001001110;
    assign rom[7'h30] = 32'b00001100000000000000000001101010;
    assign rom[7'h31] = 32'b10101101001001010000000000000100;
    assign rom[7'h32] = 32'b00001100000000000000000001101010;
    assign rom[7'h33] = 32'b10101101001000000000000000001100;
    assign rom[7'h34] = 32'b00000000000111101110100000000000;
    assign rom[7'h35] = 32'b10001111101111100000000000001000;
    assign rom[7'h36] = 32'b10001111101111110000000000001100;
    assign rom[7'h37] = 32'b00100011101111010000000000010000;
    assign rom[7'h38] = 32'b00000011111000000000000000001000;
    assign rom[7'h39] = 32'b00100011101111011111111111110000;
    assign rom[7'h3a] = 32'b10101111101111110000000000001100;
    assign rom[7'h3b] = 32'b10101111101111100000000000001000;
    assign rom[7'h3c] = 32'b00000000000111011111000000000000;
    assign rom[7'h3d] = 32'b00001100000000000000000001001110;
    assign rom[7'h3e] = 32'b00001100000000000000000001101010;
    assign rom[7'h3f] = 32'b10101101001000000000000000000000;
    assign rom[7'h40] = 32'b00110100000000100000000010100001;
    assign rom[7'h41] = 32'b00001100000000000000000001101010;
    assign rom[7'h42] = 32'b10101101001000100000000000000100;
    assign rom[7'h43] = 32'b00110100000000100000000000000001;
    assign rom[7'h44] = 32'b00001100000000000000000001101010;
    assign rom[7'h45] = 32'b10101101001000100000000000001000;
    assign rom[7'h46] = 32'b00001100000000000000000001101010;
    assign rom[7'h47] = 32'b10001101001000100000000000000000;
    assign rom[7'h48] = 32'b10101101001000000000000000001100;
    assign rom[7'h49] = 32'b00000000000111101110100000000000;
    assign rom[7'h4a] = 32'b10001111101111100000000000001000;
    assign rom[7'h4b] = 32'b10001111101111110000000000001100;
    assign rom[7'h4c] = 32'b00100011101111010000000000010000;
    assign rom[7'h4d] = 32'b00000011111000000000000000001000;
    assign rom[7'h4e] = 32'b00100011101111011111111111101100;
    assign rom[7'h4f] = 32'b10101111101111110000000000010000;
    assign rom[7'h50] = 32'b10101111101111100000000000001100;
    assign rom[7'h51] = 32'b10101111101001100000000000001000;
    assign rom[7'h52] = 32'b10101111101000100000000000000100;
    assign rom[7'h53] = 32'b00000000000111011111000000000000;
    assign rom[7'h54] = 32'b00001100000000000000000001101010;
    assign rom[7'h55] = 32'b10101101001000000000000000000000;
    assign rom[7'h56] = 32'b00110100000000100000000010100000;
    assign rom[7'h57] = 32'b00001100000000000000000001101010;
    assign rom[7'h58] = 32'b10101101001000100000000000000100;
    assign rom[7'h59] = 32'b00001100000000000000000001101010;
    assign rom[7'h5a] = 32'b10001101001001100000000000000100;
    assign rom[7'h5b] = 32'b00110000110001100000000000001000;
    assign rom[7'h5c] = 32'b00010100110000001111111111111000;
    assign rom[7'h5d] = 32'b00000000000001000001001000000010;
    assign rom[7'h5e] = 32'b00110000010000100000000000001111;
    assign rom[7'h5f] = 32'b10101101001000100000000000000100;
    assign rom[7'h60] = 32'b00110000100000100000000011111111;
    assign rom[7'h61] = 32'b00001100000000000000000001101010;
    assign rom[7'h62] = 32'b10101101001000100000000000000100;
    assign rom[7'h63] = 32'b00000000000111101110100000000000;
    assign rom[7'h64] = 32'b10001111101000100000000000000100;
    assign rom[7'h65] = 32'b10001111101001100000000000001000;
    assign rom[7'h66] = 32'b10001111101111100000000000001100;
    assign rom[7'h67] = 32'b10001111101111110000000000010000;
    assign rom[7'h68] = 32'b00100011101111010000000000010100;
    assign rom[7'h69] = 32'b00000011111000000000000000001000;
    assign rom[7'h6a] = 32'b00100011101111011111111111101100;
    assign rom[7'h6b] = 32'b10101111101111110000000000010000;
    assign rom[7'h6c] = 32'b10101111101111100000000000001100;
    assign rom[7'h6d] = 32'b10101111101001100000000000001000;
    assign rom[7'h6e] = 32'b00000000000111011111000000000000;
    assign rom[7'h6f] = 32'b10001101001001100000000000000100;
    assign rom[7'h70] = 32'b00110000110001100000000000100000;
    assign rom[7'h71] = 32'b00010000110000001111111111111101;
    assign rom[7'h72] = 32'b00000000000111101110100000000000;
    assign rom[7'h73] = 32'b10001111101001100000000000001000;
    assign rom[7'h74] = 32'b10001111101111100000000000001100;
    assign rom[7'h75] = 32'b10001111101111110000000000010000;
    assign rom[7'h76] = 32'b00100011101111010000000000010100;
    assign rom[7'h77] = 32'b00000011111000000000000000001000;
    assign rom[7'h78] = 32'b00000000000000000000000000000000;
    assign rom[7'h79] = 32'b00000000000000000000000000000000;
    assign rom[7'h7a] = 32'b00000000000000000000000000000000;
    assign rom[7'h7b] = 32'b00000000000000000000000000000000;
    assign rom[7'h7c] = 32'b00000000000000000000000000000000;
    assign rom[7'h7d] = 32'b00000000000000000000000000000000;
    assign rom[7'h7e] = 32'b00000000000000000000000000000000;
    assign rom[7'h7f] = 32'b00000000000000000000000000000000;
endmodule
