module NAND2(input logic A, 
             input logic B, 
             output logic X);
  assign X = ~(A & B);
endmodule
