package adder_pkg;

parameter N_BITS = 4;

endpackage
