package counter_pkg;

parameter N_BITS = 2;

endpackage
