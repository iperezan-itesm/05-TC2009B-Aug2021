/************************************************
  The Verilog HDL code example is from the book
  Computer Principles and Design in Verilog HDL
  by Yamin Li, published by A JOHN WILEY & SONS
************************************************/
module dec5e (n,ena,e);                  // 5-32 decoder with an enable
    input   [4:0] n;                     // 5-bit number
    input         ena;                   // master enable
    output [31:0] e;                     // 32-bit enables
    assign        e = ena? decoder(n) : 32'h00000000;
    function [31:0] decoder;
        input [4:0] n;
        case (n)
            5'd00: decoder=32'h00000001; // 00000000000000000000000000000001
            5'd01: decoder=32'h00000002; // 00000000000000000000000000000010
            5'd02: decoder=32'h00000004; // 00000000000000000000000000000100
            5'd03: decoder=32'h00000008; // 00000000000000000000000000001000
            5'd04: decoder=32'h00000010; // 00000000000000000000000000010000
            5'd05: decoder=32'h00000020; // 00000000000000000000000000100000
            5'd06: decoder=32'h00000040; // 00000000000000000000000001000000
            5'd07: decoder=32'h00000080; // 00000000000000000000000010000000
            5'd08: decoder=32'h00000100; // 00000000000000000000000100000000
            5'd09: decoder=32'h00000200; // 00000000000000000000001000000000
            5'd10: decoder=32'h00000400; // 00000000000000000000010000000000
            5'd11: decoder=32'h00000800; // 00000000000000000000100000000000
            5'd12: decoder=32'h00001000; // 00000000000000000001000000000000
            5'd13: decoder=32'h00002000; // 00000000000000000010000000000000
            5'd14: decoder=32'h00004000; // 00000000000000000100000000000000
            5'd15: decoder=32'h00008000; // 00000000000000001000000000000000
            5'd16: decoder=32'h00010000; // 00000000000000010000000000000000
            5'd17: decoder=32'h00020000; // 00000000000000100000000000000000
            5'd18: decoder=32'h00040000; // 00000000000001000000000000000000
            5'd19: decoder=32'h00080000; // 00000000000010000000000000000000
            5'd20: decoder=32'h00100000; // 00000000000100000000000000000000
            5'd21: decoder=32'h00200000; // 00000000001000000000000000000000
            5'd22: decoder=32'h00400000; // 00000000010000000000000000000000
            5'd23: decoder=32'h00800000; // 00000000100000000000000000000000
            5'd24: decoder=32'h01000000; // 00000001000000000000000000000000
            5'd25: decoder=32'h02000000; // 00000010000000000000000000000000
            5'd26: decoder=32'h04000000; // 00000100000000000000000000000000
            5'd27: decoder=32'h08000000; // 00001000000000000000000000000000
            5'd28: decoder=32'h10000000; // 00010000000000000000000000000000
            5'd29: decoder=32'h20000000; // 00100000000000000000000000000000
            5'd30: decoder=32'h40000000; // 01000000000000000000000000000000
            5'd31: decoder=32'h80000000; // 10000000000000000000000000000000
        endcase
    endfunction
endmodule
