package traffic_light_pkg;
  typedef enum logic [1:0] {
    GREEN  = 2'b00,
    YELLOW = 2'b01,
    RED    = 2'b10
  } traffic_light_t;
endpackage
